module top_module( 
    input a, b,
    output cout, sum 
);



endmodule
